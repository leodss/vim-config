//---------------------------------------------------------
//$File           : 

//$Author         : Thuan Nguyen Xuan
//$Modifier       : Thuan Nguyen Xuan

//$Created Date   : 
//$Modified Date  : 
//$Project        :
//$Module         : Module_name
//$Description    :

//$Version        :
//$Id             :
//---------------------------------------------------------

module Module_name
(

);

endmodule
